`define INST_OP_WIDTH 4
`define INST_OP_ALU_R      `INST_OP_WIDTH'd0
`define INST_OP_ALU_I      `INST_OP_WIDTH'd1
`define INST_OP_LOAD       `INST_OP_WIDTH'd2
`define INST_OP_STORE      `INST_OP_WIDTH'd3
`define INST_OP_BRANCH     `INST_OP_WIDTH'd4
`define INST_OP_JAL        `INST_OP_WIDTH'd5
`define INST_OP_JALR       `INST_OP_WIDTH'd6
`define INST_OP_LUI        `INST_OP_WIDTH'd7
`define INST_OP_AUIPC      `INST_OP_WIDTH'd8
`define INST_OP_INVALID    `INST_OP_WIDTH'd9

`define DATA_SIZE_WIDTH 2
`define DATA_SIZE_BYTE `DATA_SIZE_WIDTH'd0
`define DATA_SIZE_HALF `DATA_SIZE_WIDTH'd1
`define DATA_SIZE_WORD `DATA_SIZE_WIDTH'd2

`define EXTEND_TYPE_WIDTH 1
`define ZERO_EXTEND `EXTEND_TYPE_WIDTH'd0
`define SIGN_EXTEND `EXTEND_TYPE_WIDTH'd1
